* not(A+B+C)

*PARAMETROS
.include 32nm_HP.pm

* Declarando Fontes de tensão
Vvdd vdd gnd 1

* Declaração das fontes
Va a gnd PWL (0n 0 8n 0 8.01n 1 16n 1)
Vb b gnd PWL (0n 0 4n 0 4.01n 1 8n 1 8.01n 0 12n 0 12.01n 1 16n 1)
Vc c gnd PWL (0n 0 2n 0 2.01 1 4n 1 4.01n 0 6n 0 6.01n 1 8n 1 8.01n 0 10n 0 10.01n 1 12n 1 12.01n 0 14n 0 14.01n 1 16n 1)

* Declarando o circuito

* Declarando transistores rede pull up (em sequência)
MpA vdd a n1 vdd PMOS w=140n l=32n
MpB n1 b n2 vdd PMOS w=140n l=32n
MpC n2 c s vdd PMOS w=140n l=32n

* Declarando transistores redepull down (em paralelo)
MnA s a gnd gnd NMOS w=70n l=32n
MnB s b gnd gnd NMOS w=70n l=32n
MnB s c gnd gnd NMOS w=70n l=32n

* Simulação Transiente de 20ns com passo de 0.1ns
.tran 0.1ns 20ns 

* Fim do Arquivo SPICE
.end