*not((A+B).C)
* Declaração das fontes
Va a gnd PWL (0n 0 8n 0 8.01n 1 16n 1)
Vb b gnd PWL (0n 0 4n 0 4.01n 1 8n 1 8.01n 0 12n 0 12.01n 1 16n 1)
Vc c gnd PWL (0n 0 2n 0 2.01 1 4n 1 4.01n 0 6n 0 6.01n 1 8n 1 8.01n 0 10n 0 10.01n 1 12n 1 12.01n 0 14n 0 14.01n 1 16n 1)

* Declarando o circuito

* Declarando transistores rede pull up (A e B em sequência e C em paralelo)
MpA vdd a n1 vdd PMOS w=140n l=32n
MpB n1 b s vdd PMOS w=140n l=32n
MpC vdd c s vdd PMOS w=140n l=32n

* Declarando transistores redepull down (A e B em paralelo e C em sequência)
MnA s a n2 gnd NMOS w=70n l=32n
MnB s b n2 gnd NMOS w=70n l=32n
MnB n2 c gnd gnd NMOS w=70n l=32n

* Simulação Transiente de 20ns com passo de 0.1ns
.tran 0.1ns 20ns 

* Fim do Arquivo SPICE
.end